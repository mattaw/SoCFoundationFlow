/* Test file only */
`ifndef __WAF_TEST_INCLUDE_ONLY
`define __WAF_TEST_INCLUDE_ONLY

`endif
