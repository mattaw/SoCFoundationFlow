`define INCREMENT 1
