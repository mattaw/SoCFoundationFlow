module add_one (
    input [15:0 ] a,
    output [15:0]  b
);

assign a = b + 1;


endmodule

 
