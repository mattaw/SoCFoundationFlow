`define INCREMENT2 2
