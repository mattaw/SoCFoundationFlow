/* Pointless module part of the waf test suite */

module tb (
);

logic a;

endmodule

 
