module add_one_l2_5 (
    input [15:0 ] a,
    output [15:0]  b
);

add_one a1 (
    .a(a),
    .b(b)
);

endmodule

