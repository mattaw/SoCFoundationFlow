/* Pointless module part of the waf test suite */

module src (
    input [15:0 ] a,
    output [15:0]  b
);

assign b = a + 1;


endmodule

 
